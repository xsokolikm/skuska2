module packages #()