asdfasdfasdf asdf asdf asd fasdfasd