module produkciaBE #()