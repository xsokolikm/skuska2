module package #()