asdfasdfasdf asdf asdf asd fasdfasd asdasdasdas