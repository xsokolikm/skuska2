This is what i want to add.