module produkcia #()