asdfasdfasdf asdf asdf asd fasdf asdasd asd